module xrv1_csr
#(
    parameter ITAG_WIDTH_P = 2
) (
    ////////////////////////////////////////////////////////////////////////////////
    input logic                                 clk_i,
    input logic                                 rst_i,
    ////////////////////////////////////////////////////////////////////////////////
    output logic                                csr_rdy_o,
    input logic                                 csr_req_vld_i,
    input logic [1:0]                           csr_opc_i,
    input logic [31:0]                          csr_src0_i,
    input logic [11:0]                          csr_addr_i,
    ////////////////////////////////////////////////////////////////////////////////
    output logic                                csr_done_o,
    output logic [31:0]                         csr_data_o,
    ////////////////////////////////////////////////////////////////////////////////
    input logic [ITAG_WIDTH_P-1:0]              csr_itag_i,
    output logic [ITAG_WIDTH_P-1:0]             csr_itag_o
    ////////////////////////////////////////////////////////////////////////////////
);
    ////////////////////////////////////////////////////////////////////////////////
    assign csr_rdy_o  = 1'b1;
    assign csr_done_o = csr_req_vld_i;
    assign csr_itag_o = csr_itag_i;
    ////////////////////////////////////////////////////////////////////////////////

    ////////////////////////////////////////////////////////////////////////////////
    logic [31:0] csr_w_data_r;
    logic [31:0] csr_r_data_lo;
    ////////////////////////////////////////////////////////////////////////////////
    always_comb begin
        unique case (csr_opc_i)
            XRV_CSR_WRITE: csr_w_data_r = csr_src0_i;
            XRV_CSR_SET:   csr_w_data_r = csr_src0_i | csr_r_data_lo;
            XRV_CSR_CLR:   csr_w_data_r = ~csr_src0_i & csr_r_data_lo;
            // TODO: review this part
            // added no-lint directive as crutch to satisfy verilator
            /* verilator lint_off MULTIDRIVEN */
            XRV_CSR_READ:  csr_w_data_r = csr_src0_i;
            //
        endcase
    end
    ////////////////////////////////////////////////////////////////////////////////
    logic csr_w_en_li = csr_opc_i != XRV_CSR_READ;

    ////////////////////////////////////////////////////////////////////////////////
    // CSR File
    ////////////////////////////////////////////////////////////////////////////////
    xrv1_csrf csrf (
        ////////////////////////////////////////////////////////////////////////////////
        .clk_i                  (clk_i),
        .rst_i                  (rst_i),
        ////////////////////////////////////////////////////////////////////////////////
        .csr_addr_i             (csr_addr_i),
        .csr_r_data_o           (csr_r_data_lo),
        .csr_w_en_i             (csr_w_en_li),
        .csr_w_data_i           (csr_w_data_r)
        ////////////////////////////////////////////////////////////////////////////////
    );
    ////////////////////////////////////////////////////////////////////////////////
    assign csr_data_o = csr_r_data_lo;
    ////////////////////////////////////////////////////////////////////////////////

endmodule
