`define DEFAULT_CPU_RESET_ADDRESS 'h2000

`ifndef CPU_RESET_ADDRESS
    `define CPU_RESET_ADDRESS `DEFAULT_CPU_RESET_ADDRESS
`endif
