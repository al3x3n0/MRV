import xrv1_pkg::*;

module xrv1_csrf
(
    ////////////////////////////////////////////////////////////////////////////////
    input logic                                 clk_i,
    input logic                                 rst_i,
    ////////////////////////////////////////////////////////////////////////////////
    input  logic [11:0]                         csr_addr_i,
    output logic [31:0]                         csr_r_data_o,
    input  logic                                csr_w_en_i,
    output logic [31:0]                         csr_w_data_i
    ////////////////////////////////////////////////////////////////////////////////
);
    ////////////////////////////////////////////////////////////////////////////////
    // Machine Status Register
    ////////////////////////////////////////////////////////////////////////////////
    logic [31:0]        mstatus_q, mstatus_n_r;

    ////////////////////////////////////////////////////////////////////////////////
    // Machine Trap Vector Base Address Register
    ////////////////////////////////////////////////////////////////////////////////
    logic [31:0]        mtvec_q, mtvec_n_r;

    ////////////////////////////////////////////////////////////////////////////////
    // Machine Exception Program Counter
    ////////////////////////////////////////////////////////////////////////////////
    logic [31:0]        mepc_q, mepc_n_r;

    ////////////////////////////////////////////////////////////////////////////////
    // Machine Cause Register
    ////////////////////////////////////////////////////////////////////////////////
    logic [31:0]        mcause_q, mcause_n_r;

    ////////////////////////////////////////////////////////////////////////////////
    // Machine Scratch Register
    ////////////////////////////////////////////////////////////////////////////////
    logic [31:0]        mscratch_q, msratch_n_r;

    ////////////////////////////////////////////////////////////////////////////////
    // Machine Trap Value Register
    ////////////////////////////////////////////////////////////////////////////////
    logic [31:0]        mtval_q, mtval_n_r;

    ////////////////////////////////////////////////////////////////////////////////
    // Machine cycle counter.
    ////////////////////////////////////////////////////////////////////////////////
    logic [63:0]        mcycle_q;

    ////////////////////////////////////////////////////////////////////////////////
    always_ff @(posedge clk_i) begin
        if (rst_i) begin
            mtvec_q <= 'b0;
        end
        else if (csr_w_en_i) begin
            unique case (csr_addr_i)
                XRV_CSR_MTVEC: mtvec_q <= csr_w_data_i;
                'h7b2: mscratch_q <= csr_w_data_i;
                default:;
            endcase
        end
    end
    ////////////////////////////////////////////////////////////////////////////////

    ////////////////////////////////////////////////////////////////////////////////
    always_comb begin
        unique case (csr_addr_i)
            XRV_CSR_MTVEC: csr_r_data_o = mtvec_q;
            'h7b2: csr_r_data_o = mscratch_q;
            default: csr_r_data_o = '0;
        endcase
    end
    ////////////////////////////////////////////////////////////////////////////////

endmodule
