module mrv1_rf
#(
    ////////////////////////////////////////////////////////////////////////////////
    parameter DATA_WIDTH_P = 32,
    parameter NUM_TW_P = 8,
    parameter rf_addr_width_p = 5,
    ////////////////////////////////////////////////////////////////////////////////
    parameter twid_width_lp = $clog2(NUM_TW_P),
    parameter rf_addr_width_lp = twid_width_lp + rf_addr_width_p,
    parameter rf_size_lp = (1 << rf_addr_size_width_lp)
    ////////////////////////////////////////////////////////////////////////////////
) (
    ////////////////////////////////////////////////////////////////////////////////
    input  logic                                clk_i,
    input  logic                                rst_i,
    ////////////////////////////////////////////////////////////////////////////////
    input  logic [twid_width_lp-1:0]            twid_i,
    ////////////////////////////////////////////////////////////////////////////////
    // Read port 0
    ////////////////////////////////////////////////////////////////////////////////
    input  logic [rf_addr_width_p-1:0]          rs0_addr_i,
    output logic [DATA_WIDTH_P-1:0]             rs0_data_o,
    ////////////////////////////////////////////////////////////////////////////////
    // Read port 1
    ////////////////////////////////////////////////////////////////////////////////
    input  logic [rf_addr_width_p-1:0]          rs1_addr_i,
    output logic [DATA_WIDTH_P-1:0]             rs1_data_o,
    ////////////////////////////////////////////////////////////////////////////////
    // Write port 0
    ////////////////////////////////////////////////////////////////////////////////
    input  logic [twid_width_lp-1:0]            rd_twid_i,
    input  logic                                rd_w_en_i,
    input  logic [rf_addr_width_p-1:0]          rd_addr_i,
    input  logic [DATA_WIDTH_P-1:0]             rd_data_i
    ////////////////////////////////////////////////////////////////////////////////
);
    ////////////////////////////////////////////////////////////////////////////////
    logic [rf_size_lp-1:0][DATA_WIDTH_P-1:0]    rf_mem_q;
    ////////////////////////////////////////////////////////////////////////////////
    wire [rf_addr_width_lp-1:0] rs0_addr_w = {twid_i, rs0_addr_i};
    wire [rf_addr_width_lp-1:0] rs1_addr_w = {twid_i, rs1_addr_i};
    wire [rf_addr_width_lp-1:0] rd_addr_w  = {rd_twid_i, rd_addr_i};
    ////////////////////////////////////////////////////////////////////////////////
    assign rs0_data_o = rs0_addr_i == 'b0 ? 'b0 : rf_mem_q[rs0_addr_w];
    assign rs1_data_o = rs1_addr_i == 'b0 ? 'b0 : rf_mem_q[rs1_addr_w];
    ////////////////////////////////////////////////////////////////////////////////
    always_ff @(posedge clk_i) begin
        if (rd_w_en_i) begin
            rf_mem_q[rd_addr_w] <= rd_data_i;
        end
    end
    ////////////////////////////////////////////////////////////////////////////////
endmodule