module xrv1_branch
#(
    parameter pc_width_p = 32,
    parameter data_width_p = 32,
    parameter ITAG_WIDTH_P = "inv"
) (
    ////////////////////////////////////////////////////////////////////////////////
    input logic                             b_req_i,
    output logic                            b_rdy_o,
    input logic                             b_is_branch_i,
    input logic                             b_is_jump_i,
    ////////////////////////////////////////////////////////////////////////////////
    input logic [31:0]                      next_pc_i,
    ////////////////////////////////////////////////////////////////////////////////
    output logic                            exec_b_pc_vld_o,
    output logic [31:0]                     exec_b_pc_o,
    ////////////////////////////////////////////////////////////////////////////////
    input logic                             alu_cmp_res_i,
    ////////////////////////////////////////////////////////////////////////////////
    output logic                            b_done_o,
    output logic [31:0]                     b_wb_data_o,
    ////////////////////////////////////////////////////////////////////////////////
    input logic [ITAG_WIDTH_P-1:0]          b_itag_i,
    output logic [ITAG_WIDTH_P-1:0]         b_itag_o
    ////////////////////////////////////////////////////////////////////////////////
);
    ////////////////////////////////////////////////////////////////////////////////
    assign b_rdy_o          = 1'b1;
    assign b_done_o         = b_req_i;
    assign b_itag_o         = b_itag_i;

    ////////////////////////////////////////////////////////////////////////////////
    // Conditional branch handling
    ////////////////////////////////////////////////////////////////////////////////
    assign exec_b_pc_vld_o = b_req_i & b_is_branch_i & ~alu_cmp_res_i;
    assign exec_b_pc_o = next_pc_i;
    ////////////////////////////////////////////////////////////////////////////////
    always_comb begin
        if (b_req_i & b_is_branch_i)
            $display("next_pc_i=%h taken=%d", next_pc_i, alu_cmp_res_i);
    end


    ////////////////////////////////////////////////////////////////////////////////
    // Link Register Writeback
    ////////////////////////////////////////////////////////////////////////////////
    assign b_wb_data_o = next_pc_i;
    ////////////////////////////////////////////////////////////////////////////////

endmodule

