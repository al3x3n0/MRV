// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

////////////////////////////////////////////////////////////////////////////////
// Engineer:       Sven Stucki - svstucki@student.ethz.ch                     //
//                                                                            //
// Additional contributions by:                                               //
//                 Michael Gautschi - gautschi@iis.ee.ethz.ch                 //
//                                                                            //
// Design Name:    Compressed instruction decoder                             //
// Project Name:   RI5CY                                                      //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    Decodes RISC-V compressed instructions into their RV32     //
//                 equivalent. This module is fully combinatorial.            //
//                 Float extensions added                                     //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

import xrv1_pkg::*;

module xrv_rv16_expander
#(
    parameter fpu_en_p = 0
)
(
    ////////////////////////////////////////////////////////////////////////////////
    input  logic [31:0]         insn_i,
    output logic [31:0]         insn_o,
    output logic                illegal_insn_o
    ////////////////////////////////////////////////////////////////////////////////
);
    ////////////////////////////////////////////////////////////////////////////////
    generate
    ////////////////////////////////////////////////////////////////////////////////
    always_comb begin
        illegal_insn_o = 1'b0;
        insn_o         = '0;
        ////////////////////////////////////////////////////////////////////////////////
        unique case (insn_i[1:0])
        ////////////////////////////////////////////////////////////////////////////////
        // C0
        ////////////////////////////////////////////////////////////////////////////////
        2'b00: begin
            unique case (insn_i[15:13])
                ////////////////////////////////////////////////////////////////////////////////
                3'b000: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.addi4spn -> addi rd', x2, imm
                    ////////////////////////////////////////////////////////////////////////////////
                    insn_o = {
                        2'b0,
                        insn_i[10:7],
                        insn_i[12:11],
                        insn_i[5],
                        insn_i[6],
                        2'b00,
                        5'h02,
                        3'b000,
                        2'b01,
                        insn_i[4:2],
                        XRV_ARITH_IMM,
                        2'b11
                    };
                    if (insn_i[12:5] == 8'b0)
                        illegal_insn_o = 1'b1;
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b001: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.fld -> fld rd', imm(rs1')
                    ////////////////////////////////////////////////////////////////////////////////
                    if (fpu_en_p == 1) // insn_i[12:10]-> offset[5:3],  insn_i[6:5]-> offset[7:6]
                        insn_o = {
                            4'b0,
                            insn_i[6:5],
                            insn_i[12:10],
                            3'b000,
                            2'b01,
                            insn_i[9:7],
                            3'b011,
                            2'b01,
                            insn_i[4:2],
                            XRV_LOAD_FP,
                            2'b11
                        };
                    else
                        illegal_insn_o = 1'b1;
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b010: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.lw -> lw rd', imm(rs1')
                    ////////////////////////////////////////////////////////////////////////////////
                    insn_o = {
                        5'b0,
                        insn_i[5],
                        insn_i[12:10],
                        insn_i[6],
                        2'b00,
                        2'b01,
                        insn_i[9:7],
                        3'b010,
                        2'b01,
                        insn_i[4:2],
                        XRV_LOAD,
                        2'b11
                    };
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b011: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.flw -> flw rd', imm(rs1')
                    ////////////////////////////////////////////////////////////////////////////////
                    if (fpu_en_p == 1)
                        insn_o = {
                            5'b0,
                            insn_i[5],
                            insn_i[12:10],
                            insn_i[6],
                            2'b00, 2'b01,
                            insn_i[9:7],
                            3'b010,
                            2'b01,
                            insn_i[4:2],
                            XRV_LOAD_FP,
                            2'b11
                        };
                    else
                        illegal_insn_o = 1'b1;
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b101: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.fsd -> fsd rs2', imm(rs1')
                    ////////////////////////////////////////////////////////////////////////////////
                    if (fpu_en_p == 1) // insn_i[12:10] -> offset[5:3], insn_i[6:5] -> offset[7:6]
                        insn_o = {
                            4'b0,
                            insn_i[6:5],
                            insn_i[12],
                            2'b01,
                            insn_i[4:2],
                            2'b01,
                            insn_i[9:7],
                            3'b011,
                            insn_i[11:10],
                            3'b000,
                            XRV_STORE_FP,
                            2'b11
                        };
                    else
                        illegal_insn_o = 1'b1;
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b110: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.sw -> sw rs2', imm(rs1')
                    ////////////////////////////////////////////////////////////////////////////////
                    insn_o = {
                        5'b0,
                        insn_i[5],
                        insn_i[12],
                        2'b01,
                        insn_i[4:2],
                        2'b01,
                        insn_i[9:7],
                        3'b010,
                        insn_i[11:10],
                        insn_i[6],
                        2'b00,
                        XRV_STORE,
                        2'b11
                    };
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b111: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.fsw -> fsw rs2', imm(rs1')
                    ////////////////////////////////////////////////////////////////////////////////
                    if (fpu_en_p == 1)
                        insn_o = {
                            5'b0,
                            insn_i[5],
                            insn_i[12],
                            2'b01,
                            insn_i[4:2],
                            2'b01,
                            insn_i[9:7],
                            3'b010,
                            insn_i[11:10],
                            insn_i[6],
                            2'b00,
                            XRV_STORE_FP,
                            2'b11
                        };
                    else
                        illegal_insn_o = 1'b1;
                    end
                ////////////////////////////////////////////////////////////////////////////////
                default: begin
                    illegal_insn_o = 1'b1;
                end
                ////////////////////////////////////////////////////////////////////////////////
            endcase
        end
        ////////////////////////////////////////////////////////////////////////////////
        // C1
        ////////////////////////////////////////////////////////////////////////////////
        2'b01: begin
            unique case (insn_i[15:13])
                3'b000: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.addi -> addi rd, rd, nzimm
                    // c.nop
                    ////////////////////////////////////////////////////////////////////////////////
                    insn_o = {
                        {6{insn_i[12]}},
                        insn_i[12],
                        insn_i[6:2],
                        insn_i[11:7],
                        3'b0,
                        insn_i[11:7],
                        XRV_ARITH_IMM,
                        2'b11
                    };
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b001, 3'b101: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // 001: c.jal -> jal x1, imm
                    // 101: c.j   -> jal x0, imm
                    ////////////////////////////////////////////////////////////////////////////////
                    insn_o = {
                        insn_i[12],
                        insn_i[8],
                        insn_i[10:9],
                        insn_i[6],
                        insn_i[7],
                        insn_i[2],
                        insn_i[11],
                        insn_i[5:3],
                        {9{insn_i[12]}},
                        4'b0,
                        ~insn_i[15],
                        XRV_JAL,
                        2'b11
                    };
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b010: begin
                    if (insn_i[11:7] == 5'b0) begin
                        ////////////////////////////////////////////////////////////////////////////////
                        // Hint -> addi x0, x0, nzimm
                        ////////////////////////////////////////////////////////////////////////////////
                        insn_o = {
                            {6{insn_i[12]}},
                            insn_i[12],
                            insn_i[6:2],
                            5'b0,
                            3'b0,
                            insn_i[11:7],
                            XRV_ARITH_IMM,
                            2'b11
                        };
                    end else begin
                        ////////////////////////////////////////////////////////////////////////////////
                        // c.li -> addi rd, x0, nzimm
                        ////////////////////////////////////////////////////////////////////////////////
                        insn_o = {
                            {6{insn_i[12]}},
                            insn_i[12],
                            insn_i[6:2],
                            5'b0,
                            3'b0,
                            insn_i[11:7],
                            XRV_ARITH_IMM,
                            2'b11
                        };
                    end
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b011: begin
                    if ({insn_i[12], insn_i[6:2]} == 6'b0) begin
                        illegal_insn_o = 1'b1;
                    end else begin
                        if (insn_i[11:7] == 5'h02) begin
                            ////////////////////////////////////////////////////////////////////////////////
                            // c.addi16sp -> addi x2, x2, nzimm
                            ////////////////////////////////////////////////////////////////////////////////
                            insn_o = {
                                {3{insn_i[12]}},
                                insn_i[4:3],
                                insn_i[5],
                                insn_i[2],
                                insn_i[6],
                                4'b0,
                                5'h02,
                                3'b000,
                                5'h02,
                                XRV_ARITH_IMM,
                                2'b11
                            };
                        end else if (insn_i[11:7] == 5'b0) begin
                            ////////////////////////////////////////////////////////////////////////////////
                            // Hint -> lui x0, imm
                            ////////////////////////////////////////////////////////////////////////////////
                            insn_o = {
                                {15 {insn_i[12]}},
                                insn_i[6:2],
                                insn_i[11:7],
                                XRV_LUI,
                                2'b11
                            };
                        end else begin
                        ////////////////////////////////////////////////////////////////////////////////
                        // c.lui -> lui rd, imm
                        ////////////////////////////////////////////////////////////////////////////////
                            insn_o = {
                                {15 {insn_i[12]}},
                                insn_i[6:2],
                                insn_i[11:7],
                                XRV_LUI,
                                2'b11
                            };
                        end
                    end
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b100: begin
                    unique case (insn_i[11:10])
                        ////////////////////////////////////////////////////////////////////////////////
                        2'b00,
                        2'b01: begin
                            ////////////////////////////////////////////////////////////////////////////////
                            // 00: c.srli -> srli rd, rd, shamt
                            // 01: c.srai -> srai rd, rd, shamt
                            ////////////////////////////////////////////////////////////////////////////////
                            if (insn_i[12] == 1'b1) begin
                                ////////////////////////////////////////////////////////////////////////////////
                                // Reserved for future custom extensions (insn_o don't care)
                                ////////////////////////////////////////////////////////////////////////////////
                                insn_o = {
                                    1'b0,
                                    insn_i[10],
                                    5'b0,
                                    insn_i[6:2],
                                    2'b01,
                                    insn_i[9:7],
                                    3'b101,
                                    2'b01,
                                    insn_i[9:7],
                                    XRV_ARITH_IMM,
                                    2'b11
                                };
                                illegal_insn_o = 1'b1;
                            end else begin
                                if (insn_i[6:2] == 5'b0) begin
                                    ////////////////////////////////////////////////////////////////////////////////
                                    // Hint
                                    ////////////////////////////////////////////////////////////////////////////////
                                    insn_o = {
                                        1'b0,
                                        insn_i[10],
                                        5'b0,
                                        insn_i[6:2],
                                        2'b01,
                                        insn_i[9:7],
                                        3'b101,
                                        2'b01,
                                        insn_i[9:7],
                                        XRV_ARITH_IMM,
                                        2'b11
                                    };
                                end else begin
                                    insn_o = {
                                        1'b0,
                                        insn_i[10],
                                        5'b0,
                                        insn_i[6:2],
                                        2'b01,
                                        insn_i[9:7],
                                        3'b101,
                                        2'b01,
                                        insn_i[9:7],
                                        XRV_ARITH_IMM,
                                        2'b11
                                    };
                                end
                            end
                        end
                        ////////////////////////////////////////////////////////////////////////////////
                        2'b10: begin
                            ////////////////////////////////////////////////////////////////////////////////
                            // c.andi -> andi rd, rd, imm
                            ////////////////////////////////////////////////////////////////////////////////
                            insn_o = {
                                {6{insn_i[12]}},
                                insn_i[12],
                                insn_i[6:2],
                                2'b01,
                                insn_i[9:7],
                                3'b111,
                                2'b01,
                                insn_i[9:7],
                                XRV_ARITH_IMM,
                                2'b11
                            };
                        end
                        ////////////////////////////////////////////////////////////////////////////////
                        2'b11: begin
                            unique case ({insn_i[12], insn_i[6:5]})
                                ////////////////////////////////////////////////////////////////////////////////
                                3'b000: begin
                                    ////////////////////////////////////////////////////////////////////////////////
                                    // c.sub -> sub rd', rd', rs2'
                                    ////////////////////////////////////////////////////////////////////////////////
                                    insn_o = {
                                        2'b01,
                                        5'b0,
                                        2'b01,
                                        insn_i[4:2],
                                        2'b01,
                                        insn_i[9:7],
                                        3'b000,
                                        2'b01,
                                        insn_i[9:7],
                                        XRV_ARITH,
                                        2'b11
                                    };
                                end
                                ////////////////////////////////////////////////////////////////////////////////
                                3'b001: begin
                                    ////////////////////////////////////////////////////////////////////////////////
                                    // c.xor -> xor rd', rd', rs2'
                                    ////////////////////////////////////////////////////////////////////////////////
                                    insn_o = {
                                        7'b0,
                                        2'b01,
                                        insn_i[4:2],
                                        2'b01,
                                        insn_i[9:7],
                                        3'b100,
                                        2'b01,
                                        insn_i[9:7],
                                        XRV_ARITH,
                                        2'b11
                                    };
                                end
                                ////////////////////////////////////////////////////////////////////////////////
                                3'b010: begin
                                    ////////////////////////////////////////////////////////////////////////////////
                                    // c.or  -> or  rd', rd', rs2'
                                    ////////////////////////////////////////////////////////////////////////////////
                                    insn_o = {
                                        7'b0,
                                        2'b01,
                                        insn_i[4:2],
                                        2'b01,
                                        insn_i[9:7],
                                        3'b110,
                                        2'b01,
                                        insn_i[9:7],
                                        XRV_ARITH,
                                        2'b11
                                    };
                                end
                                ////////////////////////////////////////////////////////////////////////////////
                                3'b011: begin
                                    ////////////////////////////////////////////////////////////////////////////////
                                    // c.and -> and rd', rd', rs2'
                                    ////////////////////////////////////////////////////////////////////////////////
                                    insn_o = {
                                        7'b0,
                                        2'b01,
                                        insn_i[4:2],
                                        2'b01,
                                        insn_i[9:7],
                                        3'b111,
                                        2'b01,
                                        insn_i[9:7],
                                        XRV_ARITH,
                                        2'b11
                                    };
                                end
                                ////////////////////////////////////////////////////////////////////////////////
                                3'b100, 3'b101, 3'b110, 3'b111: begin
                                    ////////////////////////////////////////////////////////////////////////////////
                                    // 100: c.subw
                                    // 101: c.addw
                                    ////////////////////////////////////////////////////////////////////////////////
                                    illegal_insn_o = 1'b1;
                                end
                            endcase
                        end
                    endcase
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b110, 3'b111: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // 0: c.beqz -> beq rs1', x0, imm
                    // 1: c.bnez -> bne rs1', x0, imm
                    ////////////////////////////////////////////////////////////////////////////////
                    insn_o = {
                        {4{insn_i[12]}},
                        insn_i[6:5],
                        insn_i[2],
                        5'b0,
                        2'b01,
                        insn_i[9:7],
                        2'b00,
                        insn_i[13],
                        insn_i[11:10],
                        insn_i[4:3],
                        insn_i[12],
                        XRV_BRANCH,
                        2'b11
                    };
                end
            endcase
        end
        ////////////////////////////////////////////////////////////////////////////////
        // C2
        ////////////////////////////////////////////////////////////////////////////////
        2'b10: begin
            unique case (insn_i[15:13])
                ////////////////////////////////////////////////////////////////////////////////
                3'b000: begin
                    if (insn_i[12] == 1'b1) begin
                        ////////////////////////////////////////////////////////////////////////////////
                        // Reserved for future extensions (insn_o don't care)
                        ////////////////////////////////////////////////////////////////////////////////
                        insn_o = {
                            7'b0,
                            insn_i[6:2],
                            insn_i[11:7],
                            3'b001,
                            insn_i[11:7],
                            XRV_ARITH_IMM,
                            2'b11
                        };
                        illegal_insn_o = 1'b1;
                    end else begin
                        if ((insn_i[6:2] == 5'b0) || (insn_i[11:7] == 5'b0)) begin
                            ////////////////////////////////////////////////////////////////////////////////
                            // Hint -> slli rd, rd, shamt
                            ////////////////////////////////////////////////////////////////////////////////
                            insn_o = {
                                7'b0,
                                insn_i[6:2],
                                insn_i[11:7],
                                3'b001,
                                insn_i[11:7],
                                XRV_ARITH_IMM,
                                2'b11
                            };
                        end else begin
                            ////////////////////////////////////////////////////////////////////////////////
                            // c.slli -> slli rd, rd, shamt
                            ////////////////////////////////////////////////////////////////////////////////
                            insn_o = {
                                7'b0,
                                insn_i[6:2],
                                insn_i[11:7],
                                3'b001,
                                insn_i[11:7],
                                XRV_ARITH_IMM,
                                2'b11
                            };
                        end
                    end
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b001: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.fldsp -> fld rd, imm(x2)
                    ////////////////////////////////////////////////////////////////////////////////
                    if (fpu_en_p == 1) // insn_i[6:5] -> offset[4:3], insn_i[4:2] -> offset[8:6], insn_i[12] -> offset[5]
                        insn_o = {
                            3'b0,
                            insn_i[4:2],
                            insn_i[12],
                            insn_i[6:5],
                            3'b000,
                            5'h02,
                            3'b011,
                            insn_i[11:7],
                            XRV_LOAD_FP,
                            2'b11
                        };
                    else
                        illegal_insn_o = 1'b1;
                    end
                ////////////////////////////////////////////////////////////////////////////////
                3'b010: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.lwsp -> lw rd, imm(x2)
                    ////////////////////////////////////////////////////////////////////////////////
                    insn_o = {
                        4'b0,
                        insn_i[3:2],
                        insn_i[12],
                        insn_i[6:4],
                        2'b00,
                        5'h02,
                        3'b010,
                        insn_i[11:7],
                        XRV_LOAD,
                        2'b11
                    };
                    if (insn_i[11:7] == 5'b0)
                        illegal_insn_o = 1'b1;
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b011: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.flwsp -> flw rd, imm(x2)
                    ////////////////////////////////////////////////////////////////////////////////
                    if (fpu_en_p == 1)
                        insn_o = {
                            4'b0,
                            insn_i[3:2],
                            insn_i[12],
                            insn_i[6:4],
                            2'b00,
                            5'h02,
                            3'b010,
                            insn_i[11:7],
                            XRV_LOAD_FP,
                            2'b11
                        };
                    else
                        illegal_insn_o = 1'b1;
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b100: begin
                    if (insn_i[12] == 1'b0) begin
                        if (insn_i[6:2] == 5'b0) begin
                            ////////////////////////////////////////////////////////////////////////////////
                            // c.jr -> jalr x0, rd/rs1, 0
                            ////////////////////////////////////////////////////////////////////////////////
                            insn_o = {
                                12'b0,
                                insn_i[11:7],
                                3'b0,
                                5'b0,
                                XRV_JALR,
                                2'b11
                            };
                            ////////////////////////////////////////////////////////////////////////////////
                            // c.jr with rs1 = 0 is reserved
                            ////////////////////////////////////////////////////////////////////////////////
                            if (insn_i[11:7] == 5'b0)
                                illegal_insn_o = 1'b1;
                        end else begin
                            if (insn_i[11:7] == 5'b0) begin
                                ////////////////////////////////////////////////////////////////////////////////
                                // Hint -> add x0, x0, rs2
                                ////////////////////////////////////////////////////////////////////////////////
                                insn_o = {
                                    7'b0,
                                    insn_i[6:2],
                                    5'b0,
                                    3'b0,
                                    insn_i[11:7],
                                    XRV_ARITH,
                                    2'b11
                                };
                            end else begin
                                ////////////////////////////////////////////////////////////////////////////////
                                // c.mv -> add rd, x0, rs2
                                ////////////////////////////////////////////////////////////////////////////////
                                insn_o = {
                                    7'b0,
                                    insn_i[6:2],
                                    5'b0,
                                    3'b0,
                                    insn_i[11:7],
                                    XRV_ARITH,
                                    2'b11
                                };
                            end
                        end
                    end else begin
                        if (insn_i[6:2] == 5'b0) begin
                            if (insn_i[11:7] == 5'b0) begin
                                ////////////////////////////////////////////////////////////////////////////////
                                // c.ebreak -> ebreak
                                ////////////////////////////////////////////////////////////////////////////////
                                insn_o = {32'h00_10_00_73};
                            end else begin
                                ////////////////////////////////////////////////////////////////////////////////
                                // c.jalr -> jalr x1, rs1, 0
                                ////////////////////////////////////////////////////////////////////////////////
                                insn_o = {
                                    12'b0,
                                    insn_i[11:7],
                                    3'b000,
                                    5'b00001,
                                    XRV_JALR,
                                    2'b11
                                };
                            end
                        end else begin
                            if (insn_i[11:7] == 5'b0) begin
                                ////////////////////////////////////////////////////////////////////////////////
                                // Hint -> add x0, x0, rs2
                                ////////////////////////////////////////////////////////////////////////////////
                                insn_o = {
                                    7'b0,
                                    insn_i[6:2],
                                    insn_i[11:7],
                                    3'b0,
                                    insn_i[11:7],
                                    XRV_ARITH,
                                    2'b11
                                };
                            end else begin
                                ////////////////////////////////////////////////////////////////////////////////
                                // c.add -> add rd, rd, rs2
                                ////////////////////////////////////////////////////////////////////////////////
                                insn_o = {
                                    7'b0,
                                    insn_i[6:2],
                                    insn_i[11:7],
                                    3'b0,
                                    insn_i[11:7],
                                    XRV_ARITH,
                                    2'b11
                                };
                            end
                        end
                    end
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b101: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.fsdsp -> fsd rs2, imm(x2)
                    ////////////////////////////////////////////////////////////////////////////////
                    if (fpu_en_p == 1) // insn_i[12:10] -> offset[5:3], insn_i[9:7] -> offset[8:6]
                        insn_o = {
                            3'b0,
                            insn_i[9:7],
                            insn_i[12],
                            insn_i[6:2],
                            5'h02,
                            3'b011,
                            insn_i[11:10],
                            3'b000,
                            XRV_STORE_FP,
                            2'b11
                        };
                    else
                        illegal_insn_o = 1'b1;
                    end
                ////////////////////////////////////////////////////////////////////////////////
                3'b110: begin
                    ////////////////////////////////////////////////////////////////////////////////
                    // c.swsp -> sw rs2, imm(x2)
                    ////////////////////////////////////////////////////////////////////////////////
                    insn_o = {
                        4'b0,
                        insn_i[8:7],
                        insn_i[12],
                        insn_i[6:2],
                        5'h02,
                        3'b010,
                        insn_i[11:9],
                        2'b00,
                        XRV_STORE,
                        2'b11
                    };
                end
                ////////////////////////////////////////////////////////////////////////////////
                3'b111: begin
                ////////////////////////////////////////////////////////////////////////////////
                // c.fswsp -> fsw rs2, imm(x2)
                ////////////////////////////////////////////////////////////////////////////////
                if (fpu_en_p == 1)
                    insn_o = {
                        4'b0,
                        insn_i[8:7],
                        insn_i[12],
                        insn_i[6:2],
                        5'h02,
                        3'b010,
                        insn_i[11:9],
                        2'b00,
                        XRV_STORE_FP,
                        2'b11
                    };
                else
                    illegal_insn_o = 1'b1;
                end
            endcase
        end
        ////////////////////////////////////////////////////////////////////////////////
        default: begin
            insn_o = insn_i;
        end
        ////////////////////////////////////////////////////////////////////////////////
        endcase
    end
    ////////////////////////////////////////////////////////////////////////////////
    endgenerate
    ////////////////////////////////////////////////////////////////////////////////
endmodule