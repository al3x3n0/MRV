`define DEFAULT_CPU_RESET_ADDRESS 'h2000
`define DEFAULT_RAM_SIZE_BITS 16

`ifndef CPU_RESET_ADDRESS
    `define CPU_RESET_ADDRESS `DEFAULT_CPU_RESET_ADDRESS
`endif

`ifndef CPU_RAM_SIZE_BITS
    `define CPU_RAM_SIZE_BITS `DEFAULT_RAM_SIZE_BITS
`endif
