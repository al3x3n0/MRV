module xrv1_sim_ram
#(
    parameter depth_p = 1 << 16,
    parameter addr_width_lp = $clog2(depth_p)
)
(
    ////////////////////////////////////////////////////////////////////////////////
    input  logic                        clk_i,
    ////////////////////////////////////////////////////////////////////////////////
    input  logic [addr_width_lp-1:0]    addr_0_i,
    output logic [31:0]                 r_data_0_o,
    ////////////////////////////////////////////////////////////////////////////////
    input  logic [addr_width_lp-1:0]    addr_1_i,
    output logic [31:0]                 r_data_1_o,
    input  logic                        w_en_1_i,
    input  logic [31:0]                 w_data_1_i,
    input  logic [3:0]                  w_be_1_i
    ////////////////////////////////////////////////////////////////////////////////
);
    ////////////////////////////////////////////////////////////////////////////////
    logic [7:0] ram [depth_p-1:0];
    ////////////////////////////////////////////////////////////////////////////////
    wire [addr_width_lp-1:0] addr_algn0_w = {addr_0_i[addr_width_lp-1:2], 2'b00};
    wire [addr_width_lp-1:0] addr_algn1_w = {addr_1_i[addr_width_lp-1:2], 2'b00};
    ////////////////////////////////////////////////////////////////////////////////
    genvar i;
    generate
        for (i = 0; i < 4; i = i + 1) begin
            always @(posedge clk_i) begin
                ////////////////////////////////////////////////////////////////////////////////
                r_data_0_o[i * 8 +: 8] <= ram[addr_algn0_w + i];
                r_data_1_o[i * 8 +: 8] <= ram[addr_algn1_w + i];
                ////////////////////////////////////////////////////////////////////////////////
                if (w_en_1_i & w_be_1_i[i]) begin
                    ram[addr_algn1_w + i] <= w_data_1_i[i * 8 +: 8];
                end
                ////////////////////////////////////////////////////////////////////////////////
            end
        end
    endgenerate
    ////////////////////////////////////////////////////////////////////////////////

    ////////////////////////////////////////////////////////////////////////////////
    function [7:0] read_u8;
        /* verilator public */
        input integer byte_addr;
        read_u8 = ram[byte_addr];
    endfunction
    ////////////////////////////////////////////////////////////////////////////////
    task write_u8;
        /* verilator public */
        input integer byte_addr;
        input [7:0] val;
        ram[byte_addr] = val;
    endtask
    ////////////////////////////////////////////////////////////////////////////////

endmodule
